
module sky130_ef_sc_hd__decap_3();
endmodule

module sky130_ef_sc_hd__decap_4();
endmodule

module sky130_ef_sc_hd__decap_12();
endmodule