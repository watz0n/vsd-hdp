//From UCB EECS-151 FPGA Lab/Project

module uart #(
    parameter CLOCK_FREQ = 125_000_000,
    parameter MIN_BDRT = 9_600,
    parameter BAUD_BITS = $clog2((CLOCK_FREQ+(MIN_BDRT/2)-1) / (MIN_BDRT/2))
) (
    input clk,
    input reset,

    input [BAUD_BITS-1:0] baud_edge,

    input [7:0] data_in,
    input data_in_valid,
    output data_in_ready,

    output [7:0] data_out,
    output data_out_valid,
    input data_out_ready,

    input serial_in,
    output serial_out
);
    reg serial_in_reg, serial_out_reg;
    wire serial_out_tx;
    assign serial_out = serial_out_reg;
    always @ (posedge clk) begin
        serial_out_reg <= reset ? 1'b1 : serial_out_tx;
        serial_in_reg <= reset ? 1'b1 : serial_in;
    end

    uart_transmitter #(
        .CLOCK_FREQ(CLOCK_FREQ),
        .MIN_BDRT(MIN_BDRT)
    ) uatransmit (
        .clk(clk),
        .reset(reset),
        .baud_edge(baud_edge),
        .data_in(data_in),
        .data_in_valid(data_in_valid),
        .data_in_ready(data_in_ready),
        .serial_out(serial_out_tx)
    );

    uart_receiver #(
        .CLOCK_FREQ(CLOCK_FREQ),
        .MIN_BDRT(MIN_BDRT)
    ) uareceive (
        .clk(clk),
        .reset(reset),
        .baud_edge(baud_edge),
        .data_out(data_out),
        .data_out_valid(data_out_valid),
        .data_out_ready(data_out_ready),
        .serial_in(serial_in_reg)
    );
    
endmodule
